//Verilog HDL for "FA24SP25Analog", "RS-Latch" "functional"


module \RS-Latch  ( Q, QN, R, S );

  input S;
  input R;
  output Q;
  output QN;
endmodule
