//Verilog HDL for "FA24SP25Analog", "DigitalLogic_SAR" "functional"


module DigitalLogic_SAR (
	input CLK,
	input CompOut
	output [7:0] CDACOut,
	output 
);

endmodule
